// Automatically generated ROM with registered output
module neg_derivative_rom #(
    parameter DATA_WIDTH = 8,
    parameter ADDR_WIDTH = $clog2(256)
)(
    input  wire                  clk,
    input  wire [ADDR_WIDTH-1:0] addr,
    output reg  [DATA_WIDTH-1:0] dout
);

reg [DATA_WIDTH-1:0] rom_data;

always @(*) begin
    case(addr)
        8'd0: rom_data = 8'hF1;
        8'd1: rom_data = 8'hDC;
        8'd2: rom_data = 8'hBC;
        8'd3: rom_data = 8'h93;
        8'd4: rom_data = 8'h80;
        8'd5: rom_data = 8'h80;
        8'd6: rom_data = 8'h80;
        8'd7: rom_data = 8'h80;
        8'd8: rom_data = 8'h00;
        8'd9: rom_data = 8'h00;
        8'd10: rom_data = 8'h00;
        8'd11: rom_data = 8'h00;
        8'd12: rom_data = 8'h00;
        8'd13: rom_data = 8'h00;
        8'd14: rom_data = 8'h00;
        8'd15: rom_data = 8'h00;
        8'd16: rom_data = 8'hE2;
        8'd17: rom_data = 8'hB8;
        8'd18: rom_data = 8'h80;
        8'd19: rom_data = 8'h80;
        8'd20: rom_data = 8'h80;
        8'd21: rom_data = 8'h80;
        8'd22: rom_data = 8'h80;
        8'd23: rom_data = 8'h80;
        8'd24: rom_data = 8'h00;
        8'd25: rom_data = 8'h00;
        8'd26: rom_data = 8'h00;
        8'd27: rom_data = 8'h00;
        8'd28: rom_data = 8'h00;
        8'd29: rom_data = 8'h00;
        8'd30: rom_data = 8'h00;
        8'd31: rom_data = 8'h00;
        8'd32: rom_data = 8'hD3;
        8'd33: rom_data = 8'h94;
        8'd34: rom_data = 8'h80;
        8'd35: rom_data = 8'h80;
        8'd36: rom_data = 8'h80;
        8'd37: rom_data = 8'h80;
        8'd38: rom_data = 8'h80;
        8'd39: rom_data = 8'h80;
        8'd40: rom_data = 8'h00;
        8'd41: rom_data = 8'h00;
        8'd42: rom_data = 8'h00;
        8'd43: rom_data = 8'h00;
        8'd44: rom_data = 8'h00;
        8'd45: rom_data = 8'h00;
        8'd46: rom_data = 8'h00;
        8'd47: rom_data = 8'h00;
        8'd48: rom_data = 8'hC4;
        8'd49: rom_data = 8'h80;
        8'd50: rom_data = 8'h80;
        8'd51: rom_data = 8'h80;
        8'd52: rom_data = 8'h80;
        8'd53: rom_data = 8'h80;
        8'd54: rom_data = 8'h80;
        8'd55: rom_data = 8'h80;
        8'd56: rom_data = 8'h00;
        8'd57: rom_data = 8'h00;
        8'd58: rom_data = 8'h00;
        8'd59: rom_data = 8'h00;
        8'd60: rom_data = 8'h00;
        8'd61: rom_data = 8'h00;
        8'd62: rom_data = 8'h00;
        8'd63: rom_data = 8'h00;
        8'd64: rom_data = 8'hB5;
        8'd65: rom_data = 8'h80;
        8'd66: rom_data = 8'h80;
        8'd67: rom_data = 8'h80;
        8'd68: rom_data = 8'h80;
        8'd69: rom_data = 8'h80;
        8'd70: rom_data = 8'h80;
        8'd71: rom_data = 8'h80;
        8'd72: rom_data = 8'h00;
        8'd73: rom_data = 8'h00;
        8'd74: rom_data = 8'h00;
        8'd75: rom_data = 8'h00;
        8'd76: rom_data = 8'h00;
        8'd77: rom_data = 8'h00;
        8'd78: rom_data = 8'h00;
        8'd79: rom_data = 8'h00;
        8'd80: rom_data = 8'hA6;
        8'd81: rom_data = 8'h80;
        8'd82: rom_data = 8'h80;
        8'd83: rom_data = 8'h80;
        8'd84: rom_data = 8'h80;
        8'd85: rom_data = 8'h80;
        8'd86: rom_data = 8'h80;
        8'd87: rom_data = 8'h80;
        8'd88: rom_data = 8'h00;
        8'd89: rom_data = 8'h00;
        8'd90: rom_data = 8'h00;
        8'd91: rom_data = 8'h00;
        8'd92: rom_data = 8'h00;
        8'd93: rom_data = 8'h00;
        8'd94: rom_data = 8'h00;
        8'd95: rom_data = 8'h00;
        8'd96: rom_data = 8'h97;
        8'd97: rom_data = 8'h80;
        8'd98: rom_data = 8'h80;
        8'd99: rom_data = 8'h80;
        8'd100: rom_data = 8'h80;
        8'd101: rom_data = 8'h80;
        8'd102: rom_data = 8'h80;
        8'd103: rom_data = 8'h80;
        8'd104: rom_data = 8'h00;
        8'd105: rom_data = 8'h00;
        8'd106: rom_data = 8'h00;
        8'd107: rom_data = 8'h00;
        8'd108: rom_data = 8'h00;
        8'd109: rom_data = 8'h00;
        8'd110: rom_data = 8'h00;
        8'd111: rom_data = 8'h00;
        8'd112: rom_data = 8'h88;
        8'd113: rom_data = 8'h80;
        8'd114: rom_data = 8'h80;
        8'd115: rom_data = 8'h80;
        8'd116: rom_data = 8'h80;
        8'd117: rom_data = 8'h80;
        8'd118: rom_data = 8'h80;
        8'd119: rom_data = 8'h80;
        8'd120: rom_data = 8'h00;
        8'd121: rom_data = 8'h00;
        8'd122: rom_data = 8'h00;
        8'd123: rom_data = 8'h00;
        8'd124: rom_data = 8'h00;
        8'd125: rom_data = 8'h00;
        8'd126: rom_data = 8'h00;
        8'd127: rom_data = 8'h00;
        8'd128: rom_data = 8'h00;
        8'd129: rom_data = 8'h00;
        8'd130: rom_data = 8'h00;
        8'd131: rom_data = 8'h00;
        8'd132: rom_data = 8'h00;
        8'd133: rom_data = 8'h00;
        8'd134: rom_data = 8'h00;
        8'd135: rom_data = 8'h00;
        8'd136: rom_data = 8'h00;
        8'd137: rom_data = 8'h00;
        8'd138: rom_data = 8'h00;
        8'd139: rom_data = 8'h00;
        8'd140: rom_data = 8'h00;
        8'd141: rom_data = 8'h00;
        8'd142: rom_data = 8'h00;
        8'd143: rom_data = 8'h00;
        8'd144: rom_data = 8'h00;
        8'd145: rom_data = 8'h00;
        8'd146: rom_data = 8'h00;
        8'd147: rom_data = 8'h00;
        8'd148: rom_data = 8'h00;
        8'd149: rom_data = 8'h00;
        8'd150: rom_data = 8'h00;
        8'd151: rom_data = 8'h00;
        8'd152: rom_data = 8'h00;
        8'd153: rom_data = 8'h00;
        8'd154: rom_data = 8'h00;
        8'd155: rom_data = 8'h00;
        8'd156: rom_data = 8'h00;
        8'd157: rom_data = 8'h00;
        8'd158: rom_data = 8'h00;
        8'd159: rom_data = 8'h00;
        8'd160: rom_data = 8'h00;
        8'd161: rom_data = 8'h00;
        8'd162: rom_data = 8'h00;
        8'd163: rom_data = 8'h00;
        8'd164: rom_data = 8'h00;
        8'd165: rom_data = 8'h00;
        8'd166: rom_data = 8'h00;
        8'd167: rom_data = 8'h00;
        8'd168: rom_data = 8'h00;
        8'd169: rom_data = 8'h00;
        8'd170: rom_data = 8'h00;
        8'd171: rom_data = 8'h00;
        8'd172: rom_data = 8'h00;
        8'd173: rom_data = 8'h00;
        8'd174: rom_data = 8'h00;
        8'd175: rom_data = 8'h00;
        8'd176: rom_data = 8'h00;
        8'd177: rom_data = 8'h00;
        8'd178: rom_data = 8'h00;
        8'd179: rom_data = 8'h00;
        8'd180: rom_data = 8'h00;
        8'd181: rom_data = 8'h00;
        8'd182: rom_data = 8'h00;
        8'd183: rom_data = 8'h00;
        8'd184: rom_data = 8'h00;
        8'd185: rom_data = 8'h00;
        8'd186: rom_data = 8'h00;
        8'd187: rom_data = 8'h00;
        8'd188: rom_data = 8'h00;
        8'd189: rom_data = 8'h00;
        8'd190: rom_data = 8'h00;
        8'd191: rom_data = 8'h00;
        8'd192: rom_data = 8'h00;
        8'd193: rom_data = 8'h00;
        8'd194: rom_data = 8'h00;
        8'd195: rom_data = 8'h00;
        8'd196: rom_data = 8'h00;
        8'd197: rom_data = 8'h00;
        8'd198: rom_data = 8'h00;
        8'd199: rom_data = 8'h00;
        8'd200: rom_data = 8'h00;
        8'd201: rom_data = 8'h00;
        8'd202: rom_data = 8'h00;
        8'd203: rom_data = 8'h00;
        8'd204: rom_data = 8'h00;
        8'd205: rom_data = 8'h00;
        8'd206: rom_data = 8'h00;
        8'd207: rom_data = 8'h00;
        8'd208: rom_data = 8'h00;
        8'd209: rom_data = 8'h00;
        8'd210: rom_data = 8'h00;
        8'd211: rom_data = 8'h00;
        8'd212: rom_data = 8'h00;
        8'd213: rom_data = 8'h00;
        8'd214: rom_data = 8'h00;
        8'd215: rom_data = 8'h00;
        8'd216: rom_data = 8'h00;
        8'd217: rom_data = 8'h00;
        8'd218: rom_data = 8'h00;
        8'd219: rom_data = 8'h00;
        8'd220: rom_data = 8'h00;
        8'd221: rom_data = 8'h00;
        8'd222: rom_data = 8'h00;
        8'd223: rom_data = 8'h00;
        8'd224: rom_data = 8'h00;
        8'd225: rom_data = 8'h00;
        8'd226: rom_data = 8'h00;
        8'd227: rom_data = 8'h00;
        8'd228: rom_data = 8'h00;
        8'd229: rom_data = 8'h00;
        8'd230: rom_data = 8'h00;
        8'd231: rom_data = 8'h00;
        8'd232: rom_data = 8'h00;
        8'd233: rom_data = 8'h00;
        8'd234: rom_data = 8'h00;
        8'd235: rom_data = 8'h00;
        8'd236: rom_data = 8'h00;
        8'd237: rom_data = 8'h00;
        8'd238: rom_data = 8'h00;
        8'd239: rom_data = 8'h00;
        8'd240: rom_data = 8'h00;
        8'd241: rom_data = 8'h00;
        8'd242: rom_data = 8'h00;
        8'd243: rom_data = 8'h00;
        8'd244: rom_data = 8'h00;
        8'd245: rom_data = 8'h00;
        8'd246: rom_data = 8'h00;
        8'd247: rom_data = 8'h00;
        8'd248: rom_data = 8'h00;
        8'd249: rom_data = 8'h00;
        8'd250: rom_data = 8'h00;
        8'd251: rom_data = 8'h00;
        8'd252: rom_data = 8'h00;
        8'd253: rom_data = 8'h00;
        8'd254: rom_data = 8'h00;
        8'd255: rom_data = 8'h00;
        default: rom_data = {DATA_WIDTH{1'b0}};
    endcase
end

always @(posedge clk) begin
    dout <= rom_data;
end

endmodule
